netcdf test_displacement {
dimensions:
	x = 20 ;
	y = 10 ;
variables:
	float x(x) ;
	float y(y) ;
	float z(y, x) ;

// global attributes:
		:Conventions = "COARDS" ;
data:

 x = 155, 165, 175, 185, 195, 205, 215, 225, 235, 245, 255, 265, 275, 285, 
    295, 305, 315, 325, 335, 345 ;

 y = -450, -350, -250, -150, -50, 50, 150, 250, 350, 450 ;

 z =
  -147.5, -142.5, -137.5, -132.5, -127.5, -122.5, -117.5, -112.5, -107.5, 
    -102.5, -97.5, -92.5, -87.5, -82.5, -77.5, -72.5, -67.5, -62.5, -57.5, 
    -52.5,
  -97.5, -92.5, -87.5, -82.5, -77.5, -72.5, -67.5, -62.5, -57.5, -52.5, 
    -47.5, -42.5, -37.5, -32.5, -27.5, -22.5, -17.5, -12.5, -7.5, -2.5,
  -47.5, -42.5, -37.5, -32.5, -27.5, -22.5, -17.5, -12.5, -7.5, -2.5, 2.5, 
    7.5, 12.5, 17.5, 22.5, 27.5, 32.5, 37.5, 42.5, 47.5,
  2.5, 7.5, 12.5, 17.5, 22.5, 27.5, 32.5, 37.5, 42.5, 47.5, 52.5, 57.5, 62.5, 
    67.5, 72.5, 77.5, 82.5, 87.5, 92.5, 97.5,
  52.5, 57.5, 62.5, 67.5, 72.5, 77.5, 82.5, 87.5, 92.5, 97.5, 102.5, 107.5, 
    112.5, 117.5, 122.5, 127.5, 132.5, 137.5, 142.5, 147.5,
  102.5, 107.5, 112.5, 117.5, 122.5, 127.5, 132.5, 137.5, 142.5, 147.5, 
    152.5, 157.5, 162.5, 167.5, 172.5, 177.5, 182.5, 187.5, 192.5, 197.5,
  152.5, 157.5, 162.5, 167.5, 172.5, 177.5, 182.5, 187.5, 192.5, 197.5, 
    202.5, 207.5, 212.5, 217.5, 222.5, 227.5, 232.5, 237.5, 242.5, 247.5,
  202.5, 207.5, 212.5, 217.5, 222.5, 227.5, 232.5, 237.5, 242.5, 247.5, 
    252.5, 257.5, 262.5, 267.5, 272.5, 277.5, 282.5, 287.5, 292.5, 297.5,
  252.5, 257.5, 262.5, 267.5, 272.5, 277.5, 282.5, 287.5, 292.5, 297.5, 
    302.5, 307.5, 312.5, 317.5, 322.5, 327.5, 332.5, 337.5, 342.5, 347.5,
  302.5, 307.5, 312.5, 317.5, 322.5, 327.5, 332.5, 337.5, 342.5, 347.5, 
    352.5, 357.5, 362.5, 367.5, 372.5, 377.5, 382.5, 387.5, 392.5, 397.5 ;
}
