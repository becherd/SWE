netcdf test_bathymetry {
dimensions:
	x = 100 ;
	y = 50 ;
variables:
	float x(x) ;
	float y(y) ;
	float z(y, x) ;

// global attributes:
		:Conventions = "COARDS" ;
data:

 x = -245, -235, -225, -215, -205, -195, -185, -175, -165, -155, -145, -135, 
    -125, -115, -105, -95, -85, -75, -65, -55, -45, -35, -25, -15, -5, 5, 15, 
    25, 35, 45, 55, 65, 75, 85, 95, 105, 115, 125, 135, 145, 155, 165, 175, 
    185, 195, 205, 215, 225, 235, 245, 255, 265, 275, 285, 295, 305, 315, 
    325, 335, 345, 355, 365, 375, 385, 395, 405, 415, 425, 435, 445, 455, 
    465, 475, 485, 495, 505, 515, 525, 535, 545, 555, 565, 575, 585, 595, 
    605, 615, 625, 635, 645, 655, 665, 675, 685, 695, 705, 715, 725, 735, 745 ;

 y = -1225, -1175, -1125, -1075, -1025, -975, -925, -875, -825, -775, -725, 
    -675, -625, -575, -525, -475, -425, -375, -325, -275, -225, -175, -125, 
    -75, -25, 25, 75, 125, 175, 225, 275, 325, 375, 425, 475, 525, 575, 625, 
    675, 725, 775, 825, 875, 925, 975, 1025, 1075, 1125, 1175, 1225 ;

 z =
  300.125, 287.875, 275.625, 263.375, 251.125, 238.875, 226.625, 214.375, 
    202.125, 189.875, 177.625, 165.375, 153.125, 140.875, 128.625, 116.375, 
    104.125, 91.875, 79.625, 67.375, 55.125, 42.875, 30.625, 18.375, 6.125, 
    -6.125, -18.375, -30.625, -42.875, -55.125, -67.375, -79.625, -91.875, 
    -104.125, -116.375, -128.625, -140.875, -153.125, -165.375, -177.625, 
    -189.875, -202.125, -214.375, -226.625, -238.875, -251.125, -263.375, 
    -275.625, -287.875, -300.125, -312.375, -324.625, -336.875, -349.125, 
    -361.375, -373.625, -385.875, -398.125, -410.375, -422.625, -434.875, 
    -447.125, -459.375, -471.625, -483.875, -496.125, -508.375, -520.625, 
    -532.875, -545.125, -557.375, -569.625, -581.875, -594.125, -606.375, 
    -618.625, -630.875, -643.125, -655.375, -667.625, -679.875, -692.125, 
    -704.375, -716.625, -728.875, -741.125, -753.375, -765.625, -777.875, 
    -790.125, -802.375, -814.625, -826.875, -839.125, -851.375, -863.625, 
    -875.875, -888.125, -900.375, -912.625,
  287.875, 276.125, 264.375, 252.625, 240.875, 229.125, 217.375, 205.625, 
    193.875, 182.125, 170.375, 158.625, 146.875, 135.125, 123.375, 111.625, 
    99.875, 88.125, 76.375, 64.625, 52.875, 41.125, 29.375, 17.625, 5.875, 
    -5.875, -17.625, -29.375, -41.125, -52.875, -64.625, -76.375, -88.125, 
    -99.875, -111.625, -123.375, -135.125, -146.875, -158.625, -170.375, 
    -182.125, -193.875, -205.625, -217.375, -229.125, -240.875, -252.625, 
    -264.375, -276.125, -287.875, -299.625, -311.375, -323.125, -334.875, 
    -346.625, -358.375, -370.125, -381.875, -393.625, -405.375, -417.125, 
    -428.875, -440.625, -452.375, -464.125, -475.875, -487.625, -499.375, 
    -511.125, -522.875, -534.625, -546.375, -558.125, -569.875, -581.625, 
    -593.375, -605.125, -616.875, -628.625, -640.375, -652.125, -663.875, 
    -675.625, -687.375, -699.125, -710.875, -722.625, -734.375, -746.125, 
    -757.875, -769.625, -781.375, -793.125, -804.875, -816.625, -828.375, 
    -840.125, -851.875, -863.625, -875.375,
  275.625, 264.375, 253.125, 241.875, 230.625, 219.375, 208.125, 196.875, 
    185.625, 174.375, 163.125, 151.875, 140.625, 129.375, 118.125, 106.875, 
    95.625, 84.375, 73.125, 61.875, 50.625, 39.375, 28.125, 16.875, 5.625, 
    -5.625, -16.875, -28.125, -39.375, -50.625, -61.875, -73.125, -84.375, 
    -95.625, -106.875, -118.125, -129.375, -140.625, -151.875, -163.125, 
    -174.375, -185.625, -196.875, -208.125, -219.375, -230.625, -241.875, 
    -253.125, -264.375, -275.625, -286.875, -298.125, -309.375, -320.625, 
    -331.875, -343.125, -354.375, -365.625, -376.875, -388.125, -399.375, 
    -410.625, -421.875, -433.125, -444.375, -455.625, -466.875, -478.125, 
    -489.375, -500.625, -511.875, -523.125, -534.375, -545.625, -556.875, 
    -568.125, -579.375, -590.625, -601.875, -613.125, -624.375, -635.625, 
    -646.875, -658.125, -669.375, -680.625, -691.875, -703.125, -714.375, 
    -725.625, -736.875, -748.125, -759.375, -770.625, -781.875, -793.125, 
    -804.375, -815.625, -826.875, -838.125,
  263.375, 252.625, 241.875, 231.125, 220.375, 209.625, 198.875, 188.125, 
    177.375, 166.625, 155.875, 145.125, 134.375, 123.625, 112.875, 102.125, 
    91.375, 80.625, 69.875, 59.125, 48.375, 37.625, 26.875, 16.125, 5.375, 
    -5.375, -16.125, -26.875, -37.625, -48.375, -59.125, -69.875, -80.625, 
    -91.375, -102.125, -112.875, -123.625, -134.375, -145.125, -155.875, 
    -166.625, -177.375, -188.125, -198.875, -209.625, -220.375, -231.125, 
    -241.875, -252.625, -263.375, -274.125, -284.875, -295.625, -306.375, 
    -317.125, -327.875, -338.625, -349.375, -360.125, -370.875, -381.625, 
    -392.375, -403.125, -413.875, -424.625, -435.375, -446.125, -456.875, 
    -467.625, -478.375, -489.125, -499.875, -510.625, -521.375, -532.125, 
    -542.875, -553.625, -564.375, -575.125, -585.875, -596.625, -607.375, 
    -618.125, -628.875, -639.625, -650.375, -661.125, -671.875, -682.625, 
    -693.375, -704.125, -714.875, -725.625, -736.375, -747.125, -757.875, 
    -768.625, -779.375, -790.125, -800.875,
  251.125, 240.875, 230.625, 220.375, 210.125, 199.875, 189.625, 179.375, 
    169.125, 158.875, 148.625, 138.375, 128.125, 117.875, 107.625, 97.375, 
    87.125, 76.875, 66.625, 56.375, 46.125, 35.875, 25.625, 15.375, 5.125, 
    -5.125, -15.375, -25.625, -35.875, -46.125, -56.375, -66.625, -76.875, 
    -87.125, -97.375, -107.625, -117.875, -128.125, -138.375, -148.625, 
    -158.875, -169.125, -179.375, -189.625, -199.875, -210.125, -220.375, 
    -230.625, -240.875, -251.125, -261.375, -271.625, -281.875, -292.125, 
    -302.375, -312.625, -322.875, -333.125, -343.375, -353.625, -363.875, 
    -374.125, -384.375, -394.625, -404.875, -415.125, -425.375, -435.625, 
    -445.875, -456.125, -466.375, -476.625, -486.875, -497.125, -507.375, 
    -517.625, -527.875, -538.125, -548.375, -558.625, -568.875, -579.125, 
    -589.375, -599.625, -609.875, -620.125, -630.375, -640.625, -650.875, 
    -661.125, -671.375, -681.625, -691.875, -702.125, -712.375, -722.625, 
    -732.875, -743.125, -753.375, -763.625,
  238.875, 229.125, 219.375, 209.625, 199.875, 190.125, 180.375, 170.625, 
    160.875, 151.125, 141.375, 131.625, 121.875, 112.125, 102.375, 92.625, 
    82.875, 73.125, 63.375, 53.625, 43.875, 34.125, 24.375, 14.625, 4.875, 
    -4.875, -14.625, -24.375, -34.125, -43.875, -53.625, -63.375, -73.125, 
    -82.875, -92.625, -102.375, -112.125, -121.875, -131.625, -141.375, 
    -151.125, -160.875, -170.625, -180.375, -190.125, -199.875, -209.625, 
    -219.375, -229.125, -238.875, -248.625, -258.375, -268.125, -277.875, 
    -287.625, -297.375, -307.125, -316.875, -326.625, -336.375, -346.125, 
    -355.875, -365.625, -375.375, -385.125, -394.875, -404.625, -414.375, 
    -424.125, -433.875, -443.625, -453.375, -463.125, -472.875, -482.625, 
    -492.375, -502.125, -511.875, -521.625, -531.375, -541.125, -550.875, 
    -560.625, -570.375, -580.125, -589.875, -599.625, -609.375, -619.125, 
    -628.875, -638.625, -648.375, -658.125, -667.875, -677.625, -687.375, 
    -697.125, -706.875, -716.625, -726.375,
  226.625, 217.375, 208.125, 198.875, 189.625, 180.375, 171.125, 161.875, 
    152.625, 143.375, 134.125, 124.875, 115.625, 106.375, 97.125, 87.875, 
    78.625, 69.375, 60.125, 50.875, 41.625, 32.375, 23.125, 13.875, 4.625, 
    -4.625, -13.875, -23.125, -32.375, -41.625, -50.875, -60.125, -69.375, 
    -78.625, -87.875, -97.125, -106.375, -115.625, -124.875, -134.125, 
    -143.375, -152.625, -161.875, -171.125, -180.375, -189.625, -198.875, 
    -208.125, -217.375, -226.625, -235.875, -245.125, -254.375, -263.625, 
    -272.875, -282.125, -291.375, -300.625, -309.875, -319.125, -328.375, 
    -337.625, -346.875, -356.125, -365.375, -374.625, -383.875, -393.125, 
    -402.375, -411.625, -420.875, -430.125, -439.375, -448.625, -457.875, 
    -467.125, -476.375, -485.625, -494.875, -504.125, -513.375, -522.625, 
    -531.875, -541.125, -550.375, -559.625, -568.875, -578.125, -587.375, 
    -596.625, -605.875, -615.125, -624.375, -633.625, -642.875, -652.125, 
    -661.375, -670.625, -679.875, -689.125,
  214.375, 205.625, 196.875, 188.125, 179.375, 170.625, 161.875, 153.125, 
    144.375, 135.625, 126.875, 118.125, 109.375, 100.625, 91.875, 83.125, 
    74.375, 65.625, 56.875, 48.125, 39.375, 30.625, 21.875, 13.125, 4.375, 
    -4.375, -13.125, -21.875, -30.625, -39.375, -48.125, -56.875, -65.625, 
    -74.375, -83.125, -91.875, -100.625, -109.375, -118.125, -126.875, 
    -135.625, -144.375, -153.125, -161.875, -170.625, -179.375, -188.125, 
    -196.875, -205.625, -214.375, -223.125, -231.875, -240.625, -249.375, 
    -258.125, -266.875, -275.625, -284.375, -293.125, -301.875, -310.625, 
    -319.375, -328.125, -336.875, -345.625, -354.375, -363.125, -371.875, 
    -380.625, -389.375, -398.125, -406.875, -415.625, -424.375, -433.125, 
    -441.875, -450.625, -459.375, -468.125, -476.875, -485.625, -494.375, 
    -503.125, -511.875, -520.625, -529.375, -538.125, -546.875, -555.625, 
    -564.375, -573.125, -581.875, -590.625, -599.375, -608.125, -616.875, 
    -625.625, -634.375, -643.125, -651.875,
  202.125, 193.875, 185.625, 177.375, 169.125, 160.875, 152.625, 144.375, 
    136.125, 127.875, 119.625, 111.375, 103.125, 94.875, 86.625, 78.375, 
    70.125, 61.875, 53.625, 45.375, 37.125, 28.875, 20.625, 12.375, 4.125, 
    -4.125, -12.375, -20.625, -28.875, -37.125, -45.375, -53.625, -61.875, 
    -70.125, -78.375, -86.625, -94.875, -103.125, -111.375, -119.625, 
    -127.875, -136.125, -144.375, -152.625, -160.875, -169.125, -177.375, 
    -185.625, -193.875, -202.125, -210.375, -218.625, -226.875, -235.125, 
    -243.375, -251.625, -259.875, -268.125, -276.375, -284.625, -292.875, 
    -301.125, -309.375, -317.625, -325.875, -334.125, -342.375, -350.625, 
    -358.875, -367.125, -375.375, -383.625, -391.875, -400.125, -408.375, 
    -416.625, -424.875, -433.125, -441.375, -449.625, -457.875, -466.125, 
    -474.375, -482.625, -490.875, -499.125, -507.375, -515.625, -523.875, 
    -532.125, -540.375, -548.625, -556.875, -565.125, -573.375, -581.625, 
    -589.875, -598.125, -606.375, -614.625,
  189.875, 182.125, 174.375, 166.625, 158.875, 151.125, 143.375, 135.625, 
    127.875, 120.125, 112.375, 104.625, 96.875, 89.125, 81.375, 73.625, 
    65.875, 58.125, 50.375, 42.625, 34.875, 27.125, 19.375, 11.625, 3.875, 
    -3.875, -11.625, -19.375, -27.125, -34.875, -42.625, -50.375, -58.125, 
    -65.875, -73.625, -81.375, -89.125, -96.875, -104.625, -112.375, 
    -120.125, -127.875, -135.625, -143.375, -151.125, -158.875, -166.625, 
    -174.375, -182.125, -189.875, -197.625, -205.375, -213.125, -220.875, 
    -228.625, -236.375, -244.125, -251.875, -259.625, -267.375, -275.125, 
    -282.875, -290.625, -298.375, -306.125, -313.875, -321.625, -329.375, 
    -337.125, -344.875, -352.625, -360.375, -368.125, -375.875, -383.625, 
    -391.375, -399.125, -406.875, -414.625, -422.375, -430.125, -437.875, 
    -445.625, -453.375, -461.125, -468.875, -476.625, -484.375, -492.125, 
    -499.875, -507.625, -515.375, -523.125, -530.875, -538.625, -546.375, 
    -554.125, -561.875, -569.625, -577.375,
  177.625, 170.375, 163.125, 155.875, 148.625, 141.375, 134.125, 126.875, 
    119.625, 112.375, 105.125, 97.875, 90.625, 83.375, 76.125, 68.875, 
    61.625, 54.375, 47.125, 39.875, 32.625, 25.375, 18.125, 10.875, 3.625, 
    -3.625, -10.875, -18.125, -25.375, -32.625, -39.875, -47.125, -54.375, 
    -61.625, -68.875, -76.125, -83.375, -90.625, -97.875, -105.125, -112.375, 
    -119.625, -126.875, -134.125, -141.375, -148.625, -155.875, -163.125, 
    -170.375, -177.625, -184.875, -192.125, -199.375, -206.625, -213.875, 
    -221.125, -228.375, -235.625, -242.875, -250.125, -257.375, -264.625, 
    -271.875, -279.125, -286.375, -293.625, -300.875, -308.125, -315.375, 
    -322.625, -329.875, -337.125, -344.375, -351.625, -358.875, -366.125, 
    -373.375, -380.625, -387.875, -395.125, -402.375, -409.625, -416.875, 
    -424.125, -431.375, -438.625, -445.875, -453.125, -460.375, -467.625, 
    -474.875, -482.125, -489.375, -496.625, -503.875, -511.125, -518.375, 
    -525.625, -532.875, -540.125,
  165.375, 158.625, 151.875, 145.125, 138.375, 131.625, 124.875, 118.125, 
    111.375, 104.625, 97.875, 91.125, 84.375, 77.625, 70.875, 64.125, 57.375, 
    50.625, 43.875, 37.125, 30.375, 23.625, 16.875, 10.125, 3.375, -3.375, 
    -10.125, -16.875, -23.625, -30.375, -37.125, -43.875, -50.625, -57.375, 
    -64.125, -70.875, -77.625, -84.375, -91.125, -97.875, -104.625, -111.375, 
    -118.125, -124.875, -131.625, -138.375, -145.125, -151.875, -158.625, 
    -165.375, -172.125, -178.875, -185.625, -192.375, -199.125, -205.875, 
    -212.625, -219.375, -226.125, -232.875, -239.625, -246.375, -253.125, 
    -259.875, -266.625, -273.375, -280.125, -286.875, -293.625, -300.375, 
    -307.125, -313.875, -320.625, -327.375, -334.125, -340.875, -347.625, 
    -354.375, -361.125, -367.875, -374.625, -381.375, -388.125, -394.875, 
    -401.625, -408.375, -415.125, -421.875, -428.625, -435.375, -442.125, 
    -448.875, -455.625, -462.375, -469.125, -475.875, -482.625, -489.375, 
    -496.125, -502.875,
  153.125, 146.875, 140.625, 134.375, 128.125, 121.875, 115.625, 109.375, 
    103.125, 96.875, 90.625, 84.375, 78.125, 71.875, 65.625, 59.375, 53.125, 
    46.875, 40.625, 34.375, 28.125, 21.875, 15.625, 9.375, 3.125, -3.125, 
    -9.375, -15.625, -21.875, -28.125, -34.375, -40.625, -46.875, -53.125, 
    -59.375, -65.625, -71.875, -78.125, -84.375, -90.625, -96.875, -103.125, 
    -109.375, -115.625, -121.875, -128.125, -134.375, -140.625, -146.875, 
    -153.125, -159.375, -165.625, -171.875, -178.125, -184.375, -190.625, 
    -196.875, -203.125, -209.375, -215.625, -221.875, -228.125, -234.375, 
    -240.625, -246.875, -253.125, -259.375, -265.625, -271.875, -278.125, 
    -284.375, -290.625, -296.875, -303.125, -309.375, -315.625, -321.875, 
    -328.125, -334.375, -340.625, -346.875, -353.125, -359.375, -365.625, 
    -371.875, -378.125, -384.375, -390.625, -396.875, -403.125, -409.375, 
    -415.625, -421.875, -428.125, -434.375, -440.625, -446.875, -453.125, 
    -459.375, -465.625,
  140.875, 135.125, 129.375, 123.625, 117.875, 112.125, 106.375, 100.625, 
    94.875, 89.125, 83.375, 77.625, 71.875, 66.125, 60.375, 54.625, 48.875, 
    43.125, 37.375, 31.625, 25.875, 20.125, 14.375, 8.625, 2.875, -2.875, 
    -8.625, -14.375, -20.125, -25.875, -31.625, -37.375, -43.125, -48.875, 
    -54.625, -60.375, -66.125, -71.875, -77.625, -83.375, -89.125, -94.875, 
    -100.625, -106.375, -112.125, -117.875, -123.625, -129.375, -135.125, 
    -140.875, -146.625, -152.375, -158.125, -163.875, -169.625, -175.375, 
    -181.125, -186.875, -192.625, -198.375, -204.125, -209.875, -215.625, 
    -221.375, -227.125, -232.875, -238.625, -244.375, -250.125, -255.875, 
    -261.625, -267.375, -273.125, -278.875, -284.625, -290.375, -296.125, 
    -301.875, -307.625, -313.375, -319.125, -324.875, -330.625, -336.375, 
    -342.125, -347.875, -353.625, -359.375, -365.125, -370.875, -376.625, 
    -382.375, -388.125, -393.875, -399.625, -405.375, -411.125, -416.875, 
    -422.625, -428.375,
  128.625, 123.375, 118.125, 112.875, 107.625, 102.375, 97.125, 91.875, 
    86.625, 81.375, 76.125, 70.875, 65.625, 60.375, 55.125, 49.875, 44.625, 
    39.375, 34.125, 28.875, 23.625, 18.375, 13.125, 7.875, 2.625, -2.625, 
    -7.875, -13.125, -18.375, -23.625, -28.875, -34.125, -39.375, -44.625, 
    -49.875, -55.125, -60.375, -65.625, -70.875, -76.125, -81.375, -86.625, 
    -91.875, -97.125, -102.375, -107.625, -112.875, -118.125, -123.375, 
    -128.625, -133.875, -139.125, -144.375, -149.625, -154.875, -160.125, 
    -165.375, -170.625, -175.875, -181.125, -186.375, -191.625, -196.875, 
    -202.125, -207.375, -212.625, -217.875, -223.125, -228.375, -233.625, 
    -238.875, -244.125, -249.375, -254.625, -259.875, -265.125, -270.375, 
    -275.625, -280.875, -286.125, -291.375, -296.625, -301.875, -307.125, 
    -312.375, -317.625, -322.875, -328.125, -333.375, -338.625, -343.875, 
    -349.125, -354.375, -359.625, -364.875, -370.125, -375.375, -380.625, 
    -385.875, -391.125,
  116.375, 111.625, 106.875, 102.125, 97.375, 92.625, 87.875, 83.125, 78.375, 
    73.625, 68.875, 64.125, 59.375, 54.625, 49.875, 45.125, 40.375, 35.625, 
    30.875, 26.125, 21.375, 16.625, 11.875, 7.125, 2.375, -2.375, -7.125, 
    -11.875, -16.625, -21.375, -26.125, -30.875, -35.625, -40.375, -45.125, 
    -49.875, -54.625, -59.375, -64.125, -68.875, -73.625, -78.375, -83.125, 
    -87.875, -92.625, -97.375, -102.125, -106.875, -111.625, -116.375, 
    -121.125, -125.875, -130.625, -135.375, -140.125, -144.875, -149.625, 
    -154.375, -159.125, -163.875, -168.625, -173.375, -178.125, -182.875, 
    -187.625, -192.375, -197.125, -201.875, -206.625, -211.375, -216.125, 
    -220.875, -225.625, -230.375, -235.125, -239.875, -244.625, -249.375, 
    -254.125, -258.875, -263.625, -268.375, -273.125, -277.875, -282.625, 
    -287.375, -292.125, -296.875, -301.625, -306.375, -311.125, -315.875, 
    -320.625, -325.375, -330.125, -334.875, -339.625, -344.375, -349.125, 
    -353.875,
  104.125, 99.875, 95.625, 91.375, 87.125, 82.875, 78.625, 74.375, 70.125, 
    65.875, 61.625, 57.375, 53.125, 48.875, 44.625, 40.375, 36.125, 31.875, 
    27.625, 23.375, 19.125, 14.875, 10.625, 6.375, 2.125, -2.125, -6.375, 
    -10.625, -14.875, -19.125, -23.375, -27.625, -31.875, -36.125, -40.375, 
    -44.625, -48.875, -53.125, -57.375, -61.625, -65.875, -70.125, -74.375, 
    -78.625, -82.875, -87.125, -91.375, -95.625, -99.875, -104.125, -108.375, 
    -112.625, -116.875, -121.125, -125.375, -129.625, -133.875, -138.125, 
    -142.375, -146.625, -150.875, -155.125, -159.375, -163.625, -167.875, 
    -172.125, -176.375, -180.625, -184.875, -189.125, -193.375, -197.625, 
    -201.875, -206.125, -210.375, -214.625, -218.875, -223.125, -227.375, 
    -231.625, -235.875, -240.125, -244.375, -248.625, -252.875, -257.125, 
    -261.375, -265.625, -269.875, -274.125, -278.375, -282.625, -286.875, 
    -291.125, -295.375, -299.625, -303.875, -308.125, -312.375, -316.625,
  91.875, 88.125, 84.375, 80.625, 76.875, 73.125, 69.375, 65.625, 61.875, 
    58.125, 54.375, 50.625, 46.875, 43.125, 39.375, 35.625, 31.875, 28.125, 
    24.375, 20.625, 16.875, 13.125, 9.375, 5.625, 1.875, -1.875, -5.625, 
    -9.375, -13.125, -16.875, -20.625, -24.375, -28.125, -31.875, -35.625, 
    -39.375, -43.125, -46.875, -50.625, -54.375, -58.125, -61.875, -65.625, 
    -69.375, -73.125, -76.875, -80.625, -84.375, -88.125, -91.875, -95.625, 
    -99.375, -103.125, -106.875, -110.625, -114.375, -118.125, -121.875, 
    -125.625, -129.375, -133.125, -136.875, -140.625, -144.375, -148.125, 
    -151.875, -155.625, -159.375, -163.125, -166.875, -170.625, -174.375, 
    -178.125, -181.875, -185.625, -189.375, -193.125, -196.875, -200.625, 
    -204.375, -208.125, -211.875, -215.625, -219.375, -223.125, -226.875, 
    -230.625, -234.375, -238.125, -241.875, -245.625, -249.375, -253.125, 
    -256.875, -260.625, -264.375, -268.125, -271.875, -275.625, -279.375,
  79.625, 76.375, 73.125, 69.875, 66.625, 63.375, 60.125, 56.875, 53.625, 
    50.375, 47.125, 43.875, 40.625, 37.375, 34.125, 30.875, 27.625, 24.375, 
    21.125, 17.875, 14.625, 11.375, 8.125, 4.875, 1.625, -1.625, -4.875, 
    -8.125, -11.375, -14.625, -17.875, -21.125, -24.375, -27.625, -30.875, 
    -34.125, -37.375, -40.625, -43.875, -47.125, -50.375, -53.625, -56.875, 
    -60.125, -63.375, -66.625, -69.875, -73.125, -76.375, -79.625, -82.875, 
    -86.125, -89.375, -92.625, -95.875, -99.125, -102.375, -105.625, 
    -108.875, -112.125, -115.375, -118.625, -121.875, -125.125, -128.375, 
    -131.625, -134.875, -138.125, -141.375, -144.625, -147.875, -151.125, 
    -154.375, -157.625, -160.875, -164.125, -167.375, -170.625, -173.875, 
    -177.125, -180.375, -183.625, -186.875, -190.125, -193.375, -196.625, 
    -199.875, -203.125, -206.375, -209.625, -212.875, -216.125, -219.375, 
    -222.625, -225.875, -229.125, -232.375, -235.625, -238.875, -242.125,
  67.375, 64.625, 61.875, 59.125, 56.375, 53.625, 50.875, 48.125, 45.375, 
    42.625, 39.875, 37.125, 34.375, 31.625, 28.875, 26.125, 23.375, 20.625, 
    17.875, 15.125, 12.375, 9.625, 6.875, 4.125, 1.375, -1.375, -4.125, 
    -6.875, -9.625, -12.375, -15.125, -17.875, -20.625, -23.375, -26.125, 
    -28.875, -31.625, -34.375, -37.125, -39.875, -42.625, -45.375, -48.125, 
    -50.875, -53.625, -56.375, -59.125, -61.875, -64.625, -67.375, -70.125, 
    -72.875, -75.625, -78.375, -81.125, -83.875, -86.625, -89.375, -92.125, 
    -94.875, -97.625, -100.375, -103.125, -105.875, -108.625, -111.375, 
    -114.125, -116.875, -119.625, -122.375, -125.125, -127.875, -130.625, 
    -133.375, -136.125, -138.875, -141.625, -144.375, -147.125, -149.875, 
    -152.625, -155.375, -158.125, -160.875, -163.625, -166.375, -169.125, 
    -171.875, -174.625, -177.375, -180.125, -182.875, -185.625, -188.375, 
    -191.125, -193.875, -196.625, -199.375, -202.125, -204.875,
  55.125, 52.875, 50.625, 48.375, 46.125, 43.875, 41.625, 39.375, 37.125, 
    34.875, 32.625, 30.375, 28.125, 25.875, 23.625, 21.375, 19.125, 16.875, 
    14.625, 12.375, 10.125, 7.875, 5.625, 3.375, 1.125, -1.125, -3.375, 
    -5.625, -7.875, -10.125, -12.375, -14.625, -16.875, -19.125, -21.375, 
    -23.625, -25.875, -28.125, -30.375, -32.625, -34.875, -37.125, -39.375, 
    -41.625, -43.875, -46.125, -48.375, -50.625, -52.875, -55.125, -57.375, 
    -59.625, -61.875, -64.125, -66.375, -68.625, -70.875, -73.125, -75.375, 
    -77.625, -79.875, -82.125, -84.375, -86.625, -88.875, -91.125, -93.375, 
    -95.625, -97.875, -100.125, -102.375, -104.625, -106.875, -109.125, 
    -111.375, -113.625, -115.875, -118.125, -120.375, -122.625, -124.875, 
    -127.125, -129.375, -131.625, -133.875, -136.125, -138.375, -140.625, 
    -142.875, -145.125, -147.375, -149.625, -151.875, -154.125, -156.375, 
    -158.625, -160.875, -163.125, -165.375, -167.625,
  42.875, 41.125, 39.375, 37.625, 35.875, 34.125, 32.375, 30.625, 28.875, 
    27.125, 25.375, 23.625, 21.875, 20.125, 18.375, 16.625, 14.875, 13.125, 
    11.375, 9.625, 7.875, 6.125, 4.375, 2.625, 0.875, -0.875, -2.625, -4.375, 
    -6.125, -7.875, -9.625, -11.375, -13.125, -14.875, -16.625, -18.375, 
    -20.125, -21.875, -23.625, -25.375, -27.125, -28.875, -30.625, -32.375, 
    -34.125, -35.875, -37.625, -39.375, -41.125, -42.875, -44.625, -46.375, 
    -48.125, -49.875, -51.625, -53.375, -55.125, -56.875, -58.625, -60.375, 
    -62.125, -63.875, -65.625, -67.375, -69.125, -70.875, -72.625, -74.375, 
    -76.125, -77.875, -79.625, -81.375, -83.125, -84.875, -86.625, -88.375, 
    -90.125, -91.875, -93.625, -95.375, -97.125, -98.875, -100.625, -102.375, 
    -104.125, -105.875, -107.625, -109.375, -111.125, -112.875, -114.625, 
    -116.375, -118.125, -119.875, -121.625, -123.375, -125.125, -126.875, 
    -128.625, -130.375,
  30.625, 29.375, 28.125, 26.875, 25.625, 24.375, 23.125, 21.875, 20.625, 
    19.375, 18.125, 16.875, 15.625, 14.375, 13.125, 11.875, 10.625, 9.375, 
    8.125, 6.875, 5.625, 4.375, 3.125, 1.875, 0.625, -0.625, -1.875, -3.125, 
    -4.375, -5.625, -6.875, -8.125, -9.375, -10.625, -11.875, -13.125, 
    -14.375, -15.625, -16.875, -18.125, -19.375, -20.625, -21.875, -23.125, 
    -24.375, -25.625, -26.875, -28.125, -29.375, -30.625, -31.875, -33.125, 
    -34.375, -35.625, -36.875, -38.125, -39.375, -40.625, -41.875, -43.125, 
    -44.375, -45.625, -46.875, -48.125, -49.375, -50.625, -51.875, -53.125, 
    -54.375, -55.625, -56.875, -58.125, -59.375, -60.625, -61.875, -63.125, 
    -64.375, -65.625, -66.875, -68.125, -69.375, -70.625, -71.875, -73.125, 
    -74.375, -75.625, -76.875, -78.125, -79.375, -80.625, -81.875, -83.125, 
    -84.375, -85.625, -86.875, -88.125, -89.375, -90.625, -91.875, -93.125,
  18.375, 17.625, 16.875, 16.125, 15.375, 14.625, 13.875, 13.125, 12.375, 
    11.625, 10.875, 10.125, 9.375, 8.625, 7.875, 7.125, 6.375, 5.625, 4.875, 
    4.125, 3.375, 2.625, 1.875, 1.125, 0.375, -0.375, -1.125, -1.875, -2.625, 
    -3.375, -4.125, -4.875, -5.625, -6.375, -7.125, -7.875, -8.625, -9.375, 
    -10.125, -10.875, -11.625, -12.375, -13.125, -13.875, -14.625, -15.375, 
    -16.125, -16.875, -17.625, -18.375, -19.125, -19.875, -20.625, -21.375, 
    -22.125, -22.875, -23.625, -24.375, -25.125, -25.875, -26.625, -27.375, 
    -28.125, -28.875, -29.625, -30.375, -31.125, -31.875, -32.625, -33.375, 
    -34.125, -34.875, -35.625, -36.375, -37.125, -37.875, -38.625, -39.375, 
    -40.125, -40.875, -41.625, -42.375, -43.125, -43.875, -44.625, -45.375, 
    -46.125, -46.875, -47.625, -48.375, -49.125, -49.875, -50.625, -51.375, 
    -52.125, -52.875, -53.625, -54.375, -55.125, -55.875,
  6.125, 5.875, 5.625, 5.375, 5.125, 4.875, 4.625, 4.375, 4.125, 3.875, 
    3.625, 3.375, 3.125, 2.875, 2.625, 2.375, 2.125, 1.875, 1.625, 1.375, 
    1.125, 0.875, 0.625, 0.375, 0.125, -0.125, -0.375, -0.625, -0.875, 
    -1.125, -1.375, -1.625, -1.875, -2.125, -2.375, -2.625, -2.875, -3.125, 
    -3.375, -3.625, -3.875, -4.125, -4.375, -4.625, -4.875, -5.125, -5.375, 
    -5.625, -5.875, -6.125, -6.375, -6.625, -6.875, -7.125, -7.375, -7.625, 
    -7.875, -8.125, -8.375, -8.625, -8.875, -9.125, -9.375, -9.625, -9.875, 
    -10.125, -10.375, -10.625, -10.875, -11.125, -11.375, -11.625, -11.875, 
    -12.125, -12.375, -12.625, -12.875, -13.125, -13.375, -13.625, -13.875, 
    -14.125, -14.375, -14.625, -14.875, -15.125, -15.375, -15.625, -15.875, 
    -16.125, -16.375, -16.625, -16.875, -17.125, -17.375, -17.625, -17.875, 
    -18.125, -18.375, -18.625,
  -6.125, -5.875, -5.625, -5.375, -5.125, -4.875, -4.625, -4.375, -4.125, 
    -3.875, -3.625, -3.375, -3.125, -2.875, -2.625, -2.375, -2.125, -1.875, 
    -1.625, -1.375, -1.125, -0.875, -0.625, -0.375, -0.125, 0.125, 0.375, 
    0.625, 0.875, 1.125, 1.375, 1.625, 1.875, 2.125, 2.375, 2.625, 2.875, 
    3.125, 3.375, 3.625, 3.875, 4.125, 4.375, 4.625, 4.875, 5.125, 5.375, 
    5.625, 5.875, 6.125, 6.375, 6.625, 6.875, 7.125, 7.375, 7.625, 7.875, 
    8.125, 8.375, 8.625, 8.875, 9.125, 9.375, 9.625, 9.875, 10.125, 10.375, 
    10.625, 10.875, 11.125, 11.375, 11.625, 11.875, 12.125, 12.375, 12.625, 
    12.875, 13.125, 13.375, 13.625, 13.875, 14.125, 14.375, 14.625, 14.875, 
    15.125, 15.375, 15.625, 15.875, 16.125, 16.375, 16.625, 16.875, 17.125, 
    17.375, 17.625, 17.875, 18.125, 18.375, 18.625,
  -18.375, -17.625, -16.875, -16.125, -15.375, -14.625, -13.875, -13.125, 
    -12.375, -11.625, -10.875, -10.125, -9.375, -8.625, -7.875, -7.125, 
    -6.375, -5.625, -4.875, -4.125, -3.375, -2.625, -1.875, -1.125, -0.375, 
    0.375, 1.125, 1.875, 2.625, 3.375, 4.125, 4.875, 5.625, 6.375, 7.125, 
    7.875, 8.625, 9.375, 10.125, 10.875, 11.625, 12.375, 13.125, 13.875, 
    14.625, 15.375, 16.125, 16.875, 17.625, 18.375, 19.125, 19.875, 20.625, 
    21.375, 22.125, 22.875, 23.625, 24.375, 25.125, 25.875, 26.625, 27.375, 
    28.125, 28.875, 29.625, 30.375, 31.125, 31.875, 32.625, 33.375, 34.125, 
    34.875, 35.625, 36.375, 37.125, 37.875, 38.625, 39.375, 40.125, 40.875, 
    41.625, 42.375, 43.125, 43.875, 44.625, 45.375, 46.125, 46.875, 47.625, 
    48.375, 49.125, 49.875, 50.625, 51.375, 52.125, 52.875, 53.625, 54.375, 
    55.125, 55.875,
  -30.625, -29.375, -28.125, -26.875, -25.625, -24.375, -23.125, -21.875, 
    -20.625, -19.375, -18.125, -16.875, -15.625, -14.375, -13.125, -11.875, 
    -10.625, -9.375, -8.125, -6.875, -5.625, -4.375, -3.125, -1.875, -0.625, 
    0.625, 1.875, 3.125, 4.375, 5.625, 6.875, 8.125, 9.375, 10.625, 11.875, 
    13.125, 14.375, 15.625, 16.875, 18.125, 19.375, 20.625, 21.875, 23.125, 
    24.375, 25.625, 26.875, 28.125, 29.375, 30.625, 31.875, 33.125, 34.375, 
    35.625, 36.875, 38.125, 39.375, 40.625, 41.875, 43.125, 44.375, 45.625, 
    46.875, 48.125, 49.375, 50.625, 51.875, 53.125, 54.375, 55.625, 56.875, 
    58.125, 59.375, 60.625, 61.875, 63.125, 64.375, 65.625, 66.875, 68.125, 
    69.375, 70.625, 71.875, 73.125, 74.375, 75.625, 76.875, 78.125, 79.375, 
    80.625, 81.875, 83.125, 84.375, 85.625, 86.875, 88.125, 89.375, 90.625, 
    91.875, 93.125,
  -42.875, -41.125, -39.375, -37.625, -35.875, -34.125, -32.375, -30.625, 
    -28.875, -27.125, -25.375, -23.625, -21.875, -20.125, -18.375, -16.625, 
    -14.875, -13.125, -11.375, -9.625, -7.875, -6.125, -4.375, -2.625, 
    -0.875, 0.875, 2.625, 4.375, 6.125, 7.875, 9.625, 11.375, 13.125, 14.875, 
    16.625, 18.375, 20.125, 21.875, 23.625, 25.375, 27.125, 28.875, 30.625, 
    32.375, 34.125, 35.875, 37.625, 39.375, 41.125, 42.875, 44.625, 46.375, 
    48.125, 49.875, 51.625, 53.375, 55.125, 56.875, 58.625, 60.375, 62.125, 
    63.875, 65.625, 67.375, 69.125, 70.875, 72.625, 74.375, 76.125, 77.875, 
    79.625, 81.375, 83.125, 84.875, 86.625, 88.375, 90.125, 91.875, 93.625, 
    95.375, 97.125, 98.875, 100.625, 102.375, 104.125, 105.875, 107.625, 
    109.375, 111.125, 112.875, 114.625, 116.375, 118.125, 119.875, 121.625, 
    123.375, 125.125, 126.875, 128.625, 130.375,
  -55.125, -52.875, -50.625, -48.375, -46.125, -43.875, -41.625, -39.375, 
    -37.125, -34.875, -32.625, -30.375, -28.125, -25.875, -23.625, -21.375, 
    -19.125, -16.875, -14.625, -12.375, -10.125, -7.875, -5.625, -3.375, 
    -1.125, 1.125, 3.375, 5.625, 7.875, 10.125, 12.375, 14.625, 16.875, 
    19.125, 21.375, 23.625, 25.875, 28.125, 30.375, 32.625, 34.875, 37.125, 
    39.375, 41.625, 43.875, 46.125, 48.375, 50.625, 52.875, 55.125, 57.375, 
    59.625, 61.875, 64.125, 66.375, 68.625, 70.875, 73.125, 75.375, 77.625, 
    79.875, 82.125, 84.375, 86.625, 88.875, 91.125, 93.375, 95.625, 97.875, 
    100.125, 102.375, 104.625, 106.875, 109.125, 111.375, 113.625, 115.875, 
    118.125, 120.375, 122.625, 124.875, 127.125, 129.375, 131.625, 133.875, 
    136.125, 138.375, 140.625, 142.875, 145.125, 147.375, 149.625, 151.875, 
    154.125, 156.375, 158.625, 160.875, 163.125, 165.375, 167.625,
  -67.375, -64.625, -61.875, -59.125, -56.375, -53.625, -50.875, -48.125, 
    -45.375, -42.625, -39.875, -37.125, -34.375, -31.625, -28.875, -26.125, 
    -23.375, -20.625, -17.875, -15.125, -12.375, -9.625, -6.875, -4.125, 
    -1.375, 1.375, 4.125, 6.875, 9.625, 12.375, 15.125, 17.875, 20.625, 
    23.375, 26.125, 28.875, 31.625, 34.375, 37.125, 39.875, 42.625, 45.375, 
    48.125, 50.875, 53.625, 56.375, 59.125, 61.875, 64.625, 67.375, 70.125, 
    72.875, 75.625, 78.375, 81.125, 83.875, 86.625, 89.375, 92.125, 94.875, 
    97.625, 100.375, 103.125, 105.875, 108.625, 111.375, 114.125, 116.875, 
    119.625, 122.375, 125.125, 127.875, 130.625, 133.375, 136.125, 138.875, 
    141.625, 144.375, 147.125, 149.875, 152.625, 155.375, 158.125, 160.875, 
    163.625, 166.375, 169.125, 171.875, 174.625, 177.375, 180.125, 182.875, 
    185.625, 188.375, 191.125, 193.875, 196.625, 199.375, 202.125, 204.875,
  -79.625, -76.375, -73.125, -69.875, -66.625, -63.375, -60.125, -56.875, 
    -53.625, -50.375, -47.125, -43.875, -40.625, -37.375, -34.125, -30.875, 
    -27.625, -24.375, -21.125, -17.875, -14.625, -11.375, -8.125, -4.875, 
    -1.625, 1.625, 4.875, 8.125, 11.375, 14.625, 17.875, 21.125, 24.375, 
    27.625, 30.875, 34.125, 37.375, 40.625, 43.875, 47.125, 50.375, 53.625, 
    56.875, 60.125, 63.375, 66.625, 69.875, 73.125, 76.375, 79.625, 82.875, 
    86.125, 89.375, 92.625, 95.875, 99.125, 102.375, 105.625, 108.875, 
    112.125, 115.375, 118.625, 121.875, 125.125, 128.375, 131.625, 134.875, 
    138.125, 141.375, 144.625, 147.875, 151.125, 154.375, 157.625, 160.875, 
    164.125, 167.375, 170.625, 173.875, 177.125, 180.375, 183.625, 186.875, 
    190.125, 193.375, 196.625, 199.875, 203.125, 206.375, 209.625, 212.875, 
    216.125, 219.375, 222.625, 225.875, 229.125, 232.375, 235.625, 238.875, 
    242.125,
  -91.875, -88.125, -84.375, -80.625, -76.875, -73.125, -69.375, -65.625, 
    -61.875, -58.125, -54.375, -50.625, -46.875, -43.125, -39.375, -35.625, 
    -31.875, -28.125, -24.375, -20.625, -16.875, -13.125, -9.375, -5.625, 
    -1.875, 1.875, 5.625, 9.375, 13.125, 16.875, 20.625, 24.375, 28.125, 
    31.875, 35.625, 39.375, 43.125, 46.875, 50.625, 54.375, 58.125, 61.875, 
    65.625, 69.375, 73.125, 76.875, 80.625, 84.375, 88.125, 91.875, 95.625, 
    99.375, 103.125, 106.875, 110.625, 114.375, 118.125, 121.875, 125.625, 
    129.375, 133.125, 136.875, 140.625, 144.375, 148.125, 151.875, 155.625, 
    159.375, 163.125, 166.875, 170.625, 174.375, 178.125, 181.875, 185.625, 
    189.375, 193.125, 196.875, 200.625, 204.375, 208.125, 211.875, 215.625, 
    219.375, 223.125, 226.875, 230.625, 234.375, 238.125, 241.875, 245.625, 
    249.375, 253.125, 256.875, 260.625, 264.375, 268.125, 271.875, 275.625, 
    279.375,
  -104.125, -99.875, -95.625, -91.375, -87.125, -82.875, -78.625, -74.375, 
    -70.125, -65.875, -61.625, -57.375, -53.125, -48.875, -44.625, -40.375, 
    -36.125, -31.875, -27.625, -23.375, -19.125, -14.875, -10.625, -6.375, 
    -2.125, 2.125, 6.375, 10.625, 14.875, 19.125, 23.375, 27.625, 31.875, 
    36.125, 40.375, 44.625, 48.875, 53.125, 57.375, 61.625, 65.875, 70.125, 
    74.375, 78.625, 82.875, 87.125, 91.375, 95.625, 99.875, 104.125, 108.375, 
    112.625, 116.875, 121.125, 125.375, 129.625, 133.875, 138.125, 142.375, 
    146.625, 150.875, 155.125, 159.375, 163.625, 167.875, 172.125, 176.375, 
    180.625, 184.875, 189.125, 193.375, 197.625, 201.875, 206.125, 210.375, 
    214.625, 218.875, 223.125, 227.375, 231.625, 235.875, 240.125, 244.375, 
    248.625, 252.875, 257.125, 261.375, 265.625, 269.875, 274.125, 278.375, 
    282.625, 286.875, 291.125, 295.375, 299.625, 303.875, 308.125, 312.375, 
    316.625,
  -116.375, -111.625, -106.875, -102.125, -97.375, -92.625, -87.875, -83.125, 
    -78.375, -73.625, -68.875, -64.125, -59.375, -54.625, -49.875, -45.125, 
    -40.375, -35.625, -30.875, -26.125, -21.375, -16.625, -11.875, -7.125, 
    -2.375, 2.375, 7.125, 11.875, 16.625, 21.375, 26.125, 30.875, 35.625, 
    40.375, 45.125, 49.875, 54.625, 59.375, 64.125, 68.875, 73.625, 78.375, 
    83.125, 87.875, 92.625, 97.375, 102.125, 106.875, 111.625, 116.375, 
    121.125, 125.875, 130.625, 135.375, 140.125, 144.875, 149.625, 154.375, 
    159.125, 163.875, 168.625, 173.375, 178.125, 182.875, 187.625, 192.375, 
    197.125, 201.875, 206.625, 211.375, 216.125, 220.875, 225.625, 230.375, 
    235.125, 239.875, 244.625, 249.375, 254.125, 258.875, 263.625, 268.375, 
    273.125, 277.875, 282.625, 287.375, 292.125, 296.875, 301.625, 306.375, 
    311.125, 315.875, 320.625, 325.375, 330.125, 334.875, 339.625, 344.375, 
    349.125, 353.875,
  -128.625, -123.375, -118.125, -112.875, -107.625, -102.375, -97.125, 
    -91.875, -86.625, -81.375, -76.125, -70.875, -65.625, -60.375, -55.125, 
    -49.875, -44.625, -39.375, -34.125, -28.875, -23.625, -18.375, -13.125, 
    -7.875, -2.625, 2.625, 7.875, 13.125, 18.375, 23.625, 28.875, 34.125, 
    39.375, 44.625, 49.875, 55.125, 60.375, 65.625, 70.875, 76.125, 81.375, 
    86.625, 91.875, 97.125, 102.375, 107.625, 112.875, 118.125, 123.375, 
    128.625, 133.875, 139.125, 144.375, 149.625, 154.875, 160.125, 165.375, 
    170.625, 175.875, 181.125, 186.375, 191.625, 196.875, 202.125, 207.375, 
    212.625, 217.875, 223.125, 228.375, 233.625, 238.875, 244.125, 249.375, 
    254.625, 259.875, 265.125, 270.375, 275.625, 280.875, 286.125, 291.375, 
    296.625, 301.875, 307.125, 312.375, 317.625, 322.875, 328.125, 333.375, 
    338.625, 343.875, 349.125, 354.375, 359.625, 364.875, 370.125, 375.375, 
    380.625, 385.875, 391.125,
  -140.875, -135.125, -129.375, -123.625, -117.875, -112.125, -106.375, 
    -100.625, -94.875, -89.125, -83.375, -77.625, -71.875, -66.125, -60.375, 
    -54.625, -48.875, -43.125, -37.375, -31.625, -25.875, -20.125, -14.375, 
    -8.625, -2.875, 2.875, 8.625, 14.375, 20.125, 25.875, 31.625, 37.375, 
    43.125, 48.875, 54.625, 60.375, 66.125, 71.875, 77.625, 83.375, 89.125, 
    94.875, 100.625, 106.375, 112.125, 117.875, 123.625, 129.375, 135.125, 
    140.875, 146.625, 152.375, 158.125, 163.875, 169.625, 175.375, 181.125, 
    186.875, 192.625, 198.375, 204.125, 209.875, 215.625, 221.375, 227.125, 
    232.875, 238.625, 244.375, 250.125, 255.875, 261.625, 267.375, 273.125, 
    278.875, 284.625, 290.375, 296.125, 301.875, 307.625, 313.375, 319.125, 
    324.875, 330.625, 336.375, 342.125, 347.875, 353.625, 359.375, 365.125, 
    370.875, 376.625, 382.375, 388.125, 393.875, 399.625, 405.375, 411.125, 
    416.875, 422.625, 428.375,
  -153.125, -146.875, -140.625, -134.375, -128.125, -121.875, -115.625, 
    -109.375, -103.125, -96.875, -90.625, -84.375, -78.125, -71.875, -65.625, 
    -59.375, -53.125, -46.875, -40.625, -34.375, -28.125, -21.875, -15.625, 
    -9.375, -3.125, 3.125, 9.375, 15.625, 21.875, 28.125, 34.375, 40.625, 
    46.875, 53.125, 59.375, 65.625, 71.875, 78.125, 84.375, 90.625, 96.875, 
    103.125, 109.375, 115.625, 121.875, 128.125, 134.375, 140.625, 146.875, 
    153.125, 159.375, 165.625, 171.875, 178.125, 184.375, 190.625, 196.875, 
    203.125, 209.375, 215.625, 221.875, 228.125, 234.375, 240.625, 246.875, 
    253.125, 259.375, 265.625, 271.875, 278.125, 284.375, 290.625, 296.875, 
    303.125, 309.375, 315.625, 321.875, 328.125, 334.375, 340.625, 346.875, 
    353.125, 359.375, 365.625, 371.875, 378.125, 384.375, 390.625, 396.875, 
    403.125, 409.375, 415.625, 421.875, 428.125, 434.375, 440.625, 446.875, 
    453.125, 459.375, 465.625,
  -165.375, -158.625, -151.875, -145.125, -138.375, -131.625, -124.875, 
    -118.125, -111.375, -104.625, -97.875, -91.125, -84.375, -77.625, 
    -70.875, -64.125, -57.375, -50.625, -43.875, -37.125, -30.375, -23.625, 
    -16.875, -10.125, -3.375, 3.375, 10.125, 16.875, 23.625, 30.375, 37.125, 
    43.875, 50.625, 57.375, 64.125, 70.875, 77.625, 84.375, 91.125, 97.875, 
    104.625, 111.375, 118.125, 124.875, 131.625, 138.375, 145.125, 151.875, 
    158.625, 165.375, 172.125, 178.875, 185.625, 192.375, 199.125, 205.875, 
    212.625, 219.375, 226.125, 232.875, 239.625, 246.375, 253.125, 259.875, 
    266.625, 273.375, 280.125, 286.875, 293.625, 300.375, 307.125, 313.875, 
    320.625, 327.375, 334.125, 340.875, 347.625, 354.375, 361.125, 367.875, 
    374.625, 381.375, 388.125, 394.875, 401.625, 408.375, 415.125, 421.875, 
    428.625, 435.375, 442.125, 448.875, 455.625, 462.375, 469.125, 475.875, 
    482.625, 489.375, 496.125, 502.875,
  -177.625, -170.375, -163.125, -155.875, -148.625, -141.375, -134.125, 
    -126.875, -119.625, -112.375, -105.125, -97.875, -90.625, -83.375, 
    -76.125, -68.875, -61.625, -54.375, -47.125, -39.875, -32.625, -25.375, 
    -18.125, -10.875, -3.625, 3.625, 10.875, 18.125, 25.375, 32.625, 39.875, 
    47.125, 54.375, 61.625, 68.875, 76.125, 83.375, 90.625, 97.875, 105.125, 
    112.375, 119.625, 126.875, 134.125, 141.375, 148.625, 155.875, 163.125, 
    170.375, 177.625, 184.875, 192.125, 199.375, 206.625, 213.875, 221.125, 
    228.375, 235.625, 242.875, 250.125, 257.375, 264.625, 271.875, 279.125, 
    286.375, 293.625, 300.875, 308.125, 315.375, 322.625, 329.875, 337.125, 
    344.375, 351.625, 358.875, 366.125, 373.375, 380.625, 387.875, 395.125, 
    402.375, 409.625, 416.875, 424.125, 431.375, 438.625, 445.875, 453.125, 
    460.375, 467.625, 474.875, 482.125, 489.375, 496.625, 503.875, 511.125, 
    518.375, 525.625, 532.875, 540.125,
  -189.875, -182.125, -174.375, -166.625, -158.875, -151.125, -143.375, 
    -135.625, -127.875, -120.125, -112.375, -104.625, -96.875, -89.125, 
    -81.375, -73.625, -65.875, -58.125, -50.375, -42.625, -34.875, -27.125, 
    -19.375, -11.625, -3.875, 3.875, 11.625, 19.375, 27.125, 34.875, 42.625, 
    50.375, 58.125, 65.875, 73.625, 81.375, 89.125, 96.875, 104.625, 112.375, 
    120.125, 127.875, 135.625, 143.375, 151.125, 158.875, 166.625, 174.375, 
    182.125, 189.875, 197.625, 205.375, 213.125, 220.875, 228.625, 236.375, 
    244.125, 251.875, 259.625, 267.375, 275.125, 282.875, 290.625, 298.375, 
    306.125, 313.875, 321.625, 329.375, 337.125, 344.875, 352.625, 360.375, 
    368.125, 375.875, 383.625, 391.375, 399.125, 406.875, 414.625, 422.375, 
    430.125, 437.875, 445.625, 453.375, 461.125, 468.875, 476.625, 484.375, 
    492.125, 499.875, 507.625, 515.375, 523.125, 530.875, 538.625, 546.375, 
    554.125, 561.875, 569.625, 577.375,
  -202.125, -193.875, -185.625, -177.375, -169.125, -160.875, -152.625, 
    -144.375, -136.125, -127.875, -119.625, -111.375, -103.125, -94.875, 
    -86.625, -78.375, -70.125, -61.875, -53.625, -45.375, -37.125, -28.875, 
    -20.625, -12.375, -4.125, 4.125, 12.375, 20.625, 28.875, 37.125, 45.375, 
    53.625, 61.875, 70.125, 78.375, 86.625, 94.875, 103.125, 111.375, 
    119.625, 127.875, 136.125, 144.375, 152.625, 160.875, 169.125, 177.375, 
    185.625, 193.875, 202.125, 210.375, 218.625, 226.875, 235.125, 243.375, 
    251.625, 259.875, 268.125, 276.375, 284.625, 292.875, 301.125, 309.375, 
    317.625, 325.875, 334.125, 342.375, 350.625, 358.875, 367.125, 375.375, 
    383.625, 391.875, 400.125, 408.375, 416.625, 424.875, 433.125, 441.375, 
    449.625, 457.875, 466.125, 474.375, 482.625, 490.875, 499.125, 507.375, 
    515.625, 523.875, 532.125, 540.375, 548.625, 556.875, 565.125, 573.375, 
    581.625, 589.875, 598.125, 606.375, 614.625,
  -214.375, -205.625, -196.875, -188.125, -179.375, -170.625, -161.875, 
    -153.125, -144.375, -135.625, -126.875, -118.125, -109.375, -100.625, 
    -91.875, -83.125, -74.375, -65.625, -56.875, -48.125, -39.375, -30.625, 
    -21.875, -13.125, -4.375, 4.375, 13.125, 21.875, 30.625, 39.375, 48.125, 
    56.875, 65.625, 74.375, 83.125, 91.875, 100.625, 109.375, 118.125, 
    126.875, 135.625, 144.375, 153.125, 161.875, 170.625, 179.375, 188.125, 
    196.875, 205.625, 214.375, 223.125, 231.875, 240.625, 249.375, 258.125, 
    266.875, 275.625, 284.375, 293.125, 301.875, 310.625, 319.375, 328.125, 
    336.875, 345.625, 354.375, 363.125, 371.875, 380.625, 389.375, 398.125, 
    406.875, 415.625, 424.375, 433.125, 441.875, 450.625, 459.375, 468.125, 
    476.875, 485.625, 494.375, 503.125, 511.875, 520.625, 529.375, 538.125, 
    546.875, 555.625, 564.375, 573.125, 581.875, 590.625, 599.375, 608.125, 
    616.875, 625.625, 634.375, 643.125, 651.875,
  -226.625, -217.375, -208.125, -198.875, -189.625, -180.375, -171.125, 
    -161.875, -152.625, -143.375, -134.125, -124.875, -115.625, -106.375, 
    -97.125, -87.875, -78.625, -69.375, -60.125, -50.875, -41.625, -32.375, 
    -23.125, -13.875, -4.625, 4.625, 13.875, 23.125, 32.375, 41.625, 50.875, 
    60.125, 69.375, 78.625, 87.875, 97.125, 106.375, 115.625, 124.875, 
    134.125, 143.375, 152.625, 161.875, 171.125, 180.375, 189.625, 198.875, 
    208.125, 217.375, 226.625, 235.875, 245.125, 254.375, 263.625, 272.875, 
    282.125, 291.375, 300.625, 309.875, 319.125, 328.375, 337.625, 346.875, 
    356.125, 365.375, 374.625, 383.875, 393.125, 402.375, 411.625, 420.875, 
    430.125, 439.375, 448.625, 457.875, 467.125, 476.375, 485.625, 494.875, 
    504.125, 513.375, 522.625, 531.875, 541.125, 550.375, 559.625, 568.875, 
    578.125, 587.375, 596.625, 605.875, 615.125, 624.375, 633.625, 642.875, 
    652.125, 661.375, 670.625, 679.875, 689.125,
  -238.875, -229.125, -219.375, -209.625, -199.875, -190.125, -180.375, 
    -170.625, -160.875, -151.125, -141.375, -131.625, -121.875, -112.125, 
    -102.375, -92.625, -82.875, -73.125, -63.375, -53.625, -43.875, -34.125, 
    -24.375, -14.625, -4.875, 4.875, 14.625, 24.375, 34.125, 43.875, 53.625, 
    63.375, 73.125, 82.875, 92.625, 102.375, 112.125, 121.875, 131.625, 
    141.375, 151.125, 160.875, 170.625, 180.375, 190.125, 199.875, 209.625, 
    219.375, 229.125, 238.875, 248.625, 258.375, 268.125, 277.875, 287.625, 
    297.375, 307.125, 316.875, 326.625, 336.375, 346.125, 355.875, 365.625, 
    375.375, 385.125, 394.875, 404.625, 414.375, 424.125, 433.875, 443.625, 
    453.375, 463.125, 472.875, 482.625, 492.375, 502.125, 511.875, 521.625, 
    531.375, 541.125, 550.875, 560.625, 570.375, 580.125, 589.875, 599.625, 
    609.375, 619.125, 628.875, 638.625, 648.375, 658.125, 667.875, 677.625, 
    687.375, 697.125, 706.875, 716.625, 726.375,
  -251.125, -240.875, -230.625, -220.375, -210.125, -199.875, -189.625, 
    -179.375, -169.125, -158.875, -148.625, -138.375, -128.125, -117.875, 
    -107.625, -97.375, -87.125, -76.875, -66.625, -56.375, -46.125, -35.875, 
    -25.625, -15.375, -5.125, 5.125, 15.375, 25.625, 35.875, 46.125, 56.375, 
    66.625, 76.875, 87.125, 97.375, 107.625, 117.875, 128.125, 138.375, 
    148.625, 158.875, 169.125, 179.375, 189.625, 199.875, 210.125, 220.375, 
    230.625, 240.875, 251.125, 261.375, 271.625, 281.875, 292.125, 302.375, 
    312.625, 322.875, 333.125, 343.375, 353.625, 363.875, 374.125, 384.375, 
    394.625, 404.875, 415.125, 425.375, 435.625, 445.875, 456.125, 466.375, 
    476.625, 486.875, 497.125, 507.375, 517.625, 527.875, 538.125, 548.375, 
    558.625, 568.875, 579.125, 589.375, 599.625, 609.875, 620.125, 630.375, 
    640.625, 650.875, 661.125, 671.375, 681.625, 691.875, 702.125, 712.375, 
    722.625, 732.875, 743.125, 753.375, 763.625,
  -263.375, -252.625, -241.875, -231.125, -220.375, -209.625, -198.875, 
    -188.125, -177.375, -166.625, -155.875, -145.125, -134.375, -123.625, 
    -112.875, -102.125, -91.375, -80.625, -69.875, -59.125, -48.375, -37.625, 
    -26.875, -16.125, -5.375, 5.375, 16.125, 26.875, 37.625, 48.375, 59.125, 
    69.875, 80.625, 91.375, 102.125, 112.875, 123.625, 134.375, 145.125, 
    155.875, 166.625, 177.375, 188.125, 198.875, 209.625, 220.375, 231.125, 
    241.875, 252.625, 263.375, 274.125, 284.875, 295.625, 306.375, 317.125, 
    327.875, 338.625, 349.375, 360.125, 370.875, 381.625, 392.375, 403.125, 
    413.875, 424.625, 435.375, 446.125, 456.875, 467.625, 478.375, 489.125, 
    499.875, 510.625, 521.375, 532.125, 542.875, 553.625, 564.375, 575.125, 
    585.875, 596.625, 607.375, 618.125, 628.875, 639.625, 650.375, 661.125, 
    671.875, 682.625, 693.375, 704.125, 714.875, 725.625, 736.375, 747.125, 
    757.875, 768.625, 779.375, 790.125, 800.875,
  -275.625, -264.375, -253.125, -241.875, -230.625, -219.375, -208.125, 
    -196.875, -185.625, -174.375, -163.125, -151.875, -140.625, -129.375, 
    -118.125, -106.875, -95.625, -84.375, -73.125, -61.875, -50.625, -39.375, 
    -28.125, -16.875, -5.625, 5.625, 16.875, 28.125, 39.375, 50.625, 61.875, 
    73.125, 84.375, 95.625, 106.875, 118.125, 129.375, 140.625, 151.875, 
    163.125, 174.375, 185.625, 196.875, 208.125, 219.375, 230.625, 241.875, 
    253.125, 264.375, 275.625, 286.875, 298.125, 309.375, 320.625, 331.875, 
    343.125, 354.375, 365.625, 376.875, 388.125, 399.375, 410.625, 421.875, 
    433.125, 444.375, 455.625, 466.875, 478.125, 489.375, 500.625, 511.875, 
    523.125, 534.375, 545.625, 556.875, 568.125, 579.375, 590.625, 601.875, 
    613.125, 624.375, 635.625, 646.875, 658.125, 669.375, 680.625, 691.875, 
    703.125, 714.375, 725.625, 736.875, 748.125, 759.375, 770.625, 781.875, 
    793.125, 804.375, 815.625, 826.875, 838.125,
  -287.875, -276.125, -264.375, -252.625, -240.875, -229.125, -217.375, 
    -205.625, -193.875, -182.125, -170.375, -158.625, -146.875, -135.125, 
    -123.375, -111.625, -99.875, -88.125, -76.375, -64.625, -52.875, -41.125, 
    -29.375, -17.625, -5.875, 5.875, 17.625, 29.375, 41.125, 52.875, 64.625, 
    76.375, 88.125, 99.875, 111.625, 123.375, 135.125, 146.875, 158.625, 
    170.375, 182.125, 193.875, 205.625, 217.375, 229.125, 240.875, 252.625, 
    264.375, 276.125, 287.875, 299.625, 311.375, 323.125, 334.875, 346.625, 
    358.375, 370.125, 381.875, 393.625, 405.375, 417.125, 428.875, 440.625, 
    452.375, 464.125, 475.875, 487.625, 499.375, 511.125, 522.875, 534.625, 
    546.375, 558.125, 569.875, 581.625, 593.375, 605.125, 616.875, 628.625, 
    640.375, 652.125, 663.875, 675.625, 687.375, 699.125, 710.875, 722.625, 
    734.375, 746.125, 757.875, 769.625, 781.375, 793.125, 804.875, 816.625, 
    828.375, 840.125, 851.875, 863.625, 875.375,
  -300.125, -287.875, -275.625, -263.375, -251.125, -238.875, -226.625, 
    -214.375, -202.125, -189.875, -177.625, -165.375, -153.125, -140.875, 
    -128.625, -116.375, -104.125, -91.875, -79.625, -67.375, -55.125, 
    -42.875, -30.625, -18.375, -6.125, 6.125, 18.375, 30.625, 42.875, 55.125, 
    67.375, 79.625, 91.875, 104.125, 116.375, 128.625, 140.875, 153.125, 
    165.375, 177.625, 189.875, 202.125, 214.375, 226.625, 238.875, 251.125, 
    263.375, 275.625, 287.875, 300.125, 312.375, 324.625, 336.875, 349.125, 
    361.375, 373.625, 385.875, 398.125, 410.375, 422.625, 434.875, 447.125, 
    459.375, 471.625, 483.875, 496.125, 508.375, 520.625, 532.875, 545.125, 
    557.375, 569.625, 581.875, 594.125, 606.375, 618.625, 630.875, 643.125, 
    655.375, 667.625, 679.875, 692.125, 704.375, 716.625, 728.875, 741.125, 
    753.375, 765.625, 777.875, 790.125, 802.375, 814.625, 826.875, 839.125, 
    851.375, 863.625, 875.875, 888.125, 900.375, 912.625 ;
}
